`ifndef MY_IF_IN__SV
`define MY_IF_IN__SV

interface my_if_in(input clk, input rst_n);

   logic [7:0] a;
   logic [7:0] b;
   logic       valid;  
   
endinterface


`endif
